// Periodo duracion de una nota
`define T_250ms 3000000

// Divisores de la frecuencia base del 
// reloj para obtener la nota musical,
// y sus frecuencias (redondeadas)
`define FREQ_C 45977 // 261 Hz
`define FREQ_D 40955 // 293 Hz
`define FREQ_E 36474 // 329 Hz
`define FREQ_F 34383 // 349 Hz
`define FREQ_G 30612 // 391 Hz
`define FREQ_A 27272 // 440 Hz
`define FREQ_AHash 25751 // 466 Hz
`define FREQ_PlusC 22944 // 523 Hz