module main (
    // ..
);
    // ..
endmodule