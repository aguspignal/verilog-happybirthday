module main (
    // ..
);
    // ..
    // .. test
endmodule